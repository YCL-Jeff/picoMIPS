// File Name    : opcodes.sv
// Function     : picoMIPS/Southampton Lab opcode and type definitions
// Author       : tjk, ycl (modified)
// Last rev.    : April 2025

// Include guard
`ifndef OPCODES_SV
`define OPCODES_SV

// --- Opcodes (Macro Definitions) ---
`define MUL 6'b000001
`define ADD 6'b000010
`define END 6'b000011


`endif // OPCODES_SV